//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package apb_seq_pkg;

   import uvm_pkg::*;
   import spi_cfg_pkg::*;
  
   `include "uvm_macros.svh"
   `include "base_seq.sv"
   `include "rst_seq.sv"
   `include "apb_demo_seq.sv"
   `include "spi_demo_seq.sv"
   
endpackage
