//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package spi_slave_agent_pkg;
   
   import uvm_pkg::*;
   import spi_cfg_pkg::*;
   // todo:
   // import spi_tlm package here
   
   `include "uvm_macros.svh"
   `include "spi_slave_monitor.sv"
   `include "spi_slave_agent.sv"

endpackage
