//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package spi_env_pkg;

   import uvm_pkg::*;
   import apb_agent_pkg::*;
   import spi_agent_pkg::*;
   import spi_slave_agent_pkg::*;
   import apb_slave_agent_pkg::*;
   import spi_chk_pkg::*;
   
   `include "uvm_macros.svh"
   `include "spi_env.svh"
   
endpackage
