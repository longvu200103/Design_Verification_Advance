//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package apb_seq_pkg;

   import uvm_pkg::*;
   import spi_cfg_pkg::*;
  
   `include "uvm_macros.svh"
   `include "apb_demo_seq.sv"
   
endpackage
