//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package spi_cov_pkg;

   import uvm_pkg::*;
   
   `include "uvm_macros.svh"
   `include "spi_cov.sv"
   
endpackage
