//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package apb_agent_pkg;
   import uvm_pkg::*;

   `include "uvm_macros.svh"
   `include "uvm_tb_defines.sv"

endpackage

